5 5 1
141 25 0
W 3 4 9 5 141
W 4 1 9 5 141
W 4 4 9 5 138
W 4 2 12 5 137
W 1 4 9 5 124
W 4 0 9 5 112
W 3 3 9 5 110
W 2 3 9 5 110
W 1 2 9 5 109
W 3 2 9 5 109
W 2 2 9 5 108
W 4 3 9 5 108
W 2 1 9 5 107
W 2 4 9 5 106
W 0 3 9 5 106
W 1 0 9 5 106
W 3 0 9 5 105
W 1 3 9 5 104
W 2 0 9 5 103
W 0 2 9 5 103
W 3 1 9 5 102
W 0 4 9 5 102
W 0 1 9 5 101
W 1 1 9 5 99
W 0 0 9 5 98
#ZAPIS GRY WIRTUALNY SWIAT v2.0#
#Damian Jankowski s188597#
#znak polX polY sila inicjatywa wiek#
#[A]ntylopa [C]zlowiek [S]uperman [L]is [O]wca [W]ilk [Z]olw#
#[B]arszcz [G]uarana [M]lecz [T]rawa [X]Wilczejagody#
#Superman - czlowiek z wlaczona umiejetnoscia#
